LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;

ENTITY rom IS
GENERIC ( n : integer := 24);
	PORT(
		clk : IN std_logic;
		we  : IN std_logic;
		address : IN  std_logic_vector(5 DOWNTO 0);
		datain  : IN  std_logic_vector(n-1 DOWNTO 0);
		dataout : OUT std_logic_vector(n-1 DOWNTO 0));
END ENTITY rom;

ARCHITECTURE syncroma OF rom IS

	TYPE rom_type IS ARRAY(0 TO 511) OF std_logic_vector(n-1 DOWNTO 0);
	SIGNAL rom : rom_type := (
		0 => "001000101000101001000000"
		1 => "011010000000000000010000"
		2 => "010100000000000000000000"
		3 => "000000000000000000000001"
		4 => "000000000000000000000000"
		5 => "000000000000000000000000"
		6 => "000000000000000000000000"
		7 => "000000000000000000000000"
		8 => "000000000000000000000000"
		9 => "000000000000000000000000"
		10 => "000000000000000000000000"
		11 => "000000000000000000000000"
		12 => "000000000000000000000000"
		13 => "000000000000000000000000"
		14 => "000000000000000000000000"
		15 => "000000000000000000000000"
		16 => "000000000000000000000000"
		17 => "000000000000000000000000"
		18 => "000000000000000000000000"
		19 => "000000000000000000000000"
		20 => "000000000000000000000000"
		21 => "000000000000000000000000"
		22 => "000000000000000000000000"
		23 => "000000000000000000000000"
		24 => "000000000000000000000000"
		25 => "000000000000000000000000"
		26 => "000000000000000000000000"
		27 => "000000000000000000000000"
		28 => "000000000000000000000000"
		29 => "000000000000000000000000"
		30 => "000000000000000000000000"
		31 => "000000000000000000000000"
		32 => "000000000100000000000000"
		33 => "001000100000000100000000"
		34 => "011010000000000000000000"
		35 => "000000000000000000001011"
		36 => "000000000000000000000000"
		37 => "000000000000000000000000"
		38 => "000000000000000000000000"
		39 => "101000100100001100000000"
		40 => "011100110100000000000000"
		41 => "111000010000000010010000"
		42 => "101000100100001100000000"
		43 => "011100110100000000000000"
		44 => "001000110000000010010000"
		45 => "000010100100010000000000"
		46 => "011000100100010000000000"
		47 => "011110000000000000000000"
		48 => "000000000000000000001011"
		49 => "101000100100010000000000"
		50 => "011001101000000001010000"
		51 => "010010000000000000000000"
		52 => "101000100100010000000000"
		53 => "011001101000000001010000"
		54 => "010110000000000000000000"
		55 => "000000000000000000001011"
		56 => "000000000000000000000000"
		57 => "000000000000000000000000"
		58 => "000000000000000000000000"
		59 => "000000000000000000000000"
		60 => "000000000000000000000000"
		61 => "000000000000000000000000"
		62 => "000000000000000000000000"
		63 => "000000000000000000000000"
		64 => "000000000000000000000000"
		65 => "100000011000000000000000"
		66 => "000000000000000000000101"
		67 => "000000000000000000000000"
		68 => "000000000000000000000000"
		69 => "000000000000000000000000"
		70 => "000000000000000000000000"
		71 => "000000000000000000000000"
		72 => "000000000000000000000000"
		73 => "100000001000000001010000"
		74 => "000000000000000000000101"
		75 => "000000000000000000000000"
		76 => "000000000000000000000000"
		77 => "000000000000000000000000"
		78 => "000000000000000000000000"
		79 => "000000000000000000000000"
		80 => "000000000000000000000000"
		81 => "100000101000000101000000"
		82 => "011001000000000000010000"
		83 => "000000000000000000000101"
		84 => "000000000000000000000000"
		85 => "000000000000000000000000"
		86 => "000000000000000000000000"
		87 => "000000000000000000000000"
		88 => "000000000000000000000000"
		89 => "000000000000000000000000"
		90 => "000000000000000000000000"
		91 => "000000000000000000000000"
		92 => "000000000000000000000000"
		93 => "000000000000000000000000"
		94 => "000000000000000000000000"
		95 => "000000000000000000000000"
		96 => "000000000000000000000000"
		97 => "100000100000011000000000"
		98 => "011000101000000001010000"
		99 => "000000000000000000000101"
		100 => "000000000000000000000000"
		101 => "000000000000000000000000"
		102 => "000000000000000000000000"
		103 => "000000000000000000000000"
		104 => "000000000000000000000000"
		105 => "000000000000000000000000"
		106 => "000000000000000000000000"
		107 => "000000000000000000000000"
		108 => "000000000000000000000000"
		109 => "000000000000000000000000"
		110 => "000000000000000000000000"
		111 => "000000000000000000000000"
		112 => "000000000000000000000000"
		113 => "001000101000000101000000"
		114 => "011010000000000000010000"
		115 => "010000000100000000000000"
		116 => "100000100000000100000000"
		117 => "011000001000000001010000"
		118 => "000000000000000000000101"
		119 => "000000000000000000000000"
		120 => "010000001000000001010000"
		121 => "010001000000000000000000"
		122 => "000000000000000000000011"
		123 => "000000000000000000000000"
		124 => "000000000000000000000000"
		125 => "000000000000000000000000"
		126 => "000000000000000000000000"
		127 => "000000000000000000000000"
		128 => "000000000000000000000000"
		129 => "101000000100000000000000"
		130 => "000000000000000000000111"
		131 => "000000000000000000000000"
		132 => "000000000000000000000000"
		133 => "000000000000000000000000"
		134 => "000000000000000000000000"
		135 => "000000000000000000000000"
		136 => "000000000000000000000000"
		137 => "101000001000000001010000"
		138 => "000000000000000000000111"
		139 => "000000000000000000000000"
		140 => "000000000000000000000000"
		141 => "000000000000000000000000"
		142 => "000000000000000000000000"
		143 => "000000000000000000000000"
		144 => "000000000000000000000000"
		145 => "101000101000000101000000"
		146 => "011001100000000000010000"
		147 => "000000000000000000000111"
		148 => "000000000000000000000000"
		149 => "000000000000000000000000"
		150 => "000000000000000000000000"
		151 => "000000000000000000000000"
		152 => "000000000000000000000000"
		153 => "000000000000000000000000"
		154 => "000000000000000000000000"
		155 => "000000000000000000000000"
		156 => "000000000000000000000000"
		157 => "000000000000000000000000"
		158 => "000000000000000000000000"
		159 => "000000000000000000000000"
		160 => "000000000000000000000000"
		161 => "101000100000011000000000"
		162 => "011001101000000001010000"
		163 => "000000000000000000000111"
		164 => "000000000000000000000000"
		165 => "000000000000000000000000"
		166 => "000000000000000000000000"
		167 => "000000000000000000000000"
		168 => "000000000000000000000000"
		169 => "000000000000000000000000"
		170 => "000000000000000000000000"
		171 => "000000000000000000000000"
		172 => "000000000000000000000000"
		173 => "000000000000000000000000"
		174 => "000000000000000000000000"
		175 => "000000000000000000000000"
		176 => "000000000000000000000000"
		177 => "001000101000000101000000"
		178 => "011010000000000000010000"
		179 => "010000000100000000000000"
		180 => "101000100000000100000000"
		181 => "011000001000000001010000"
		182 => "000000000000000000000111"
		183 => "000000000000000000000000"
		184 => "010000001000000001010000"
		185 => "010000000100000000000000"
		186 => "000000000000000000001001"
		187 => "000000000000000000000000"
		188 => "000000000000000000000000"
		189 => "000000000000000000000000"
		190 => "000000000000000000000000"
		191 => "000000000000000000000000"
		192 => "000000000000000000000000"
		193 => "000000000000000000000000"
		194 => "000000000000000000000000"
		195 => "000000000000000000000000"
		196 => "000000000000000000000000"
		197 => "000000000000000000000000"
		198 => "000000000000000000000000"
		199 => "000000000000000000000000"
		200 => "000000000000000000000000"
		201 => "000000000000000000000000"
		202 => "000000000000000000000000"
		203 => "000000000000000000000000"
		204 => "000000000000000000000000"
		205 => "000000000000000000000000"
		206 => "000000000000000000000000"
		207 => "000000000000000000000000"
		208 => "000000000000000000000000"
		209 => "001000101001010001000000"
		210 => "011010000000000000000000"
		211 => "100000100001010100000000"
		212 => "011001000000000000010000"
		213 => "010000000100000000000000"
		214 => "100000001000000000000000"
		215 => "001000010000000010000000"
		216 => "000000100010000000000000"
		217 => "011010000000000000010000"
		218 => "000000000000000000001011"
		219 => "100000001000000001010000"
		220 => "010010000000000000000000"
		221 => "000000000000000000001011"
		222 => "000000000000000000000000"
		223 => "000000000000000000000000"
		224 => "000000000000000000000000"
		225 => "000000000000000000000000"
		226 => "000000000000000000000000"
		227 => "000000000000000000000000"
		228 => "000000000000000000000000"
		229 => "000000000000000000000000"
		230 => "000000000000000000000000"
		231 => "000000000000000000000000"
		232 => "000000000000000000000000"
		233 => "000000000000000000000000"
		234 => "000000000000000000000000"
		235 => "000000000000000000000000"
		236 => "000000000000000000000000"
		237 => "000000000000000000000000"
		238 => "000000000000000000000000"
		239 => "000000000000000000000000"
		240 => "000000000000000000000000"
		241 => "000000000000000000000000"
		242 => "000000000000000000000000"
		243 => "000000000000000000000000"
		244 => "000000000000000000000000"
		245 => "000000000000000000000000"
		246 => "000000000000000000000000"
		247 => "000000000000000000000000"
		248 => "000000000000000000000000"
		249 => "000000000000000000000000"
		250 => "000000000000000000000000"
		251 => "000000000000000000000000"
		252 => "000000000000000000000000"
		253 => "000000000000000000000000"
		254 => "000000000000000000000000"
		255 => "000000000000000000000000"
		256 => "000000000000000000000000"
		257 => "000000000000000000000000"
		258 => "000000000000000000000000"
		259 => "000000000000000000000000"
		260 => "000000000000000000000000"
		261 => "000000000000000000000000"
		262 => "000000000000000000000000"
		263 => "000000000000000000000000"
		264 => "000000000000000000000000"
		265 => "000000000000000000000000"
		266 => "000000000000000000000000"
		267 => "000000000000000000000000"
		268 => "000000000000000000000000"
		269 => "000000000000000000000000"
		270 => "000000000000000000000000"
		271 => "000000000000000000000000"
		272 => "000000000000000000000000"
		273 => "000000000000000000000000"
		274 => "000000000000000000000000"
		275 => "000000000000000000000000"
		276 => "000000000000000000000000"
		277 => "000000000000000000000000"
		278 => "000000000000000000000000"
		279 => "000000000000000000000000"
		280 => "000000000000000000000000"
		281 => "000000000000000000000000"
		282 => "000000000000000000000000"
		283 => "000000000000000000000000"
		284 => "000000000000000000000000"
		285 => "000000000000000000000000"
		286 => "000000000000000000000000"
		287 => "000000000000000000000000"
		288 => "000000000000000000000000"
		289 => "000000000000000000000000"
		290 => "000000000000000000000000"
		291 => "000000000000000000000000"
		292 => "000000000000000000000000"
		293 => "000000000000000000000000"
		294 => "000000000000000000000000"
		295 => "000000000000000000000000"
		296 => "000000000000000000000000"
		297 => "000000000000000000000000"
		298 => "000000000000000000000000"
		299 => "000000000000000000000000"
		300 => "000000000000000000000000"
		301 => "000000000000000000000000"
		302 => "000000000000000000000000"
		303 => "000000000000000000000000"
		304 => "000000000000000000000000"
		305 => "000000000000000000000000"
		306 => "000000000000000000000000"
		307 => "000000000000000000000000"
		308 => "000000000000000000000000"
		309 => "000000000000000000000000"
		310 => "000000000000000000000000"
		311 => "000000000000000000000000"
		312 => "110000100001001100000000"
		313 => "000000000000000000001001"
		314 => "110000100010000100000000"
		315 => "000000000000000000001001"
		316 => "110000100010010100000000"
		317 => "000000000000000000001001"
		318 => "110000100010011000000000"
		319 => "000000000000000000001001"
		320 => "110000100010001000000000"
		321 => "000000000000000000001001"
		322 => "110000100010100000000000"
		323 => "000000000000000000001001"
		324 => "110000100010100100000000"
		325 => "000000000000000000001001"
		326 => "110000100010101000000000"
		327 => "000000000000000000001001"
		328 => "110000100011011000000000"
		329 => "000000000000000000001001"
		330 => "000000100010010000000000"
		331 => "000000000000000000001001"
		332 => "000000100010001100000000"
		333 => "000000000000000000001001"
		334 => "000000100000011100000000"
		335 => "000000000000000000001001"
		336 => "000000100010101100000000"
		337 => "000000000000000000001001"
		338 => "000000100010110000000000"
		339 => "000000000000000000001001"
		340 => "000000100010110100000000"
		341 => "000000000000000000001001"
		342 => "000000100010111100000000"
		343 => "000000000000000000001001"
		344 => "000000100011000000000000"
		345 => "000000000000000000001001"
		346 => "000000100011000100000000"
		347 => "000000000000000000001001"
		348 => "000000000000000000000000"
		349 => "000000000000000000000000"
		350 => "000000000000000000000000"
		351 => "000000000000000000000000"
		352 => "000000000000000000000000"
		353 => "000000000000000000000000"
		354 => "000000000000000000000000"
		355 => "000000000000000000000000"
		356 => "000000000000000000000000"
		357 => "011001100000000000000000"
		358 => "000000000000000000001011"
		359 => "011000010000000010010000"
		360 => "000000000000000000001011"
		OTHERS => X"FFFFFFFF"
		) ;
	
	BEGIN
		PROCESS(clk) IS
			BEGIN
				IF rising_edge(clk) THEN  
					IF we = '1' THEN
						rom(to_integer(unsigned(address))) <= datain;
					END IF;
				END IF;
		END PROCESS;
		dataout <= rom(to_integer(unsigned(address)));
END syncroma;